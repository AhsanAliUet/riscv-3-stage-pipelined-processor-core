/////////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2022 UET Lahore (All Rights Reserved)
//
// Project Name: RISC-V Core
// Module Name:  [forwarding_unit]
// Designer:     [AHSAN ALI]
// Description:  [The unit to solve RAW data hazards in RISC-V Core]
//
/////////////////////////////////////////////////////////////////////////////////

module forwarding_unit
   import riscv_pkg::var;
# (
   parameter  PARAM1 = VAL1,
   parameter  PARAM1 = VAL1
) (
   input  logic       clk_i,
   input  logic       rst_i,
   input  logic [3:0] input_1,
   input  logic       input_2,
   input  logic       input_3,
   output logic [3:0] output_1,
);

/////////////////////////////////////////////////////////////////////////////////
   // Local Parameters

/////////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////////////
   // Functions

/////////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////////////
   // Signals

/////////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////////////
   // Assignments and Instantiations

/////////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////////////
   // Always Statements

/////////////////////////////////////////////////////////////////////////////////

endmodule: forwarding_unit