
module encoder_2x1 #(
    parameter W = 1
)(
    input  logic in0,
    input  logic in1,

    output logic out,
);




endmodule